package pkgs;
`include "uvm_macros.svh"
import uvm_pkg::*;

`include "xtn.sv"
`include "config.sv"
//`include "interface.sv"
`include "driver.sv"
`include "driver2.sv"
`include "driver3.sv"
`include "driver4.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "sequencer.sv"
`include "sequencer2.sv"
`include "sequencer3.sv"
`include "sequencer4.sv"
`include "agent.sv"
`include "agent2.sv"
`include "Agent3.sv"
`include "agent4.sv"
`include "sequence.sv"
`include "env.sv"
`include "test.sv"

endpackage
